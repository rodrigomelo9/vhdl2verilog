module types ();

   reg signed [31:0] int_r, int_a, int_b;
   reg        [31:0] nat_r, nat_a, nat_b;
   reg        [31:0] pos_r, pos_a, pos_b;
   reg signed  [7:0] sig_r, sig_a, sig_b;
   reg         [7:0] uns_r, uns_a, uns_b;

   initial begin
      $display("Integer");
      int_a = 9;
      int_b = 2;
      int_r = int_a + int_b; $display("%1d",int_r);
      int_r = int_a - int_b; $display("%1d",int_r);
      int_r = int_a * int_b; $display("%1d",int_r);
      int_r = int_a / int_b; $display("%1d",int_r);
      int_a = 9;
      int_b = -2;
      int_r = int_a + int_b; $display("%1d",int_r);
      int_r = int_a - int_b; $display("%1d",int_r);
      int_r = int_a * int_b; $display("%1d",int_r);
      int_r = int_a / int_b; $display("%1d",int_r);
      int_a = -9;
      int_b = 2;
      int_r = int_a + int_b; $display("%1d",int_r);
      int_r = int_a - int_b; $display("%1d",int_r);
      int_r = int_a * int_b; $display("%1d",int_r);
      int_r = int_a / int_b; $display("%1d",int_r);
      int_a = -9;
      int_b = -2;
      int_r = int_a + int_b; $display("%1d",int_r);
      int_r = int_a - int_b; $display("%1d",int_r);
      int_r = int_a * int_b; $display("%1d",int_r);
      int_r = int_a / int_b; $display("%1d",int_r);
      int_r = -int_r;        $display("%1d",int_r);
      $display("Natural");
      nat_a = 9;
      nat_b = 2;
      nat_r = nat_a + nat_b; $display("%1d",nat_r);
      nat_r = nat_a - nat_b; $display("%1d",nat_r);
      nat_r = nat_a * nat_b; $display("%1d",nat_r);
      nat_r = nat_a / nat_b; $display("%1d",nat_r);
      $display("Positive");
      pos_a = 9;
      pos_b = 2;
      pos_r = pos_a + pos_b; $display("%1d",pos_r);
      pos_r = pos_a - pos_b; $display("%1d",pos_r);
      pos_r = pos_a * pos_b; $display("%1d",pos_r);
      pos_r = pos_a / pos_b; $display("%1d",pos_r);
      $display("Signed");
      sig_a = 9;
      sig_b = 2;
      sig_r = sig_a + sig_b; $display("%1d",sig_r);
      sig_r = sig_a - sig_b; $display("%1d",sig_r);
      sig_r = sig_a * sig_b; $display("%1d",sig_r);
      sig_r = sig_a / sig_b; $display("%1d",sig_r);
      sig_a = 9;
      sig_b = -2;
      sig_r = sig_a + sig_b; $display("%1d",sig_r);
      sig_r = sig_a - sig_b; $display("%1d",sig_r);
      sig_r = sig_a * sig_b; $display("%1d",sig_r);
      sig_r = sig_a / sig_b; $display("%1d",sig_r);
      sig_a = -9;
      sig_b = 2;
      sig_r = sig_a + sig_b; $display("%1d",sig_r);
      sig_r = sig_a - sig_b; $display("%1d",sig_r);
      sig_r = sig_a * sig_b; $display("%1d",sig_r);
      sig_r = sig_a / sig_b; $display("%1d",sig_r);
      sig_a = -9;
      sig_b = -2;
      sig_r = sig_a + sig_b; $display("%1d",sig_r);
      sig_r = sig_a - sig_b; $display("%1d",sig_r);
      sig_r = sig_a * sig_b; $display("%1d",sig_r);
      sig_r = sig_a / sig_b; $display("%1d",sig_r);
      sig_r = -sig_r;        $display("%1d",sig_r);
      $display("Unsigned");
      uns_a = 9;
      uns_b = 2;
      uns_r = uns_a + uns_b; $display("%1d",uns_r);
      uns_r = uns_a - uns_b; $display("%1d",uns_r);
      uns_r = uns_a * uns_b; $display("%1d",uns_r);
      uns_r = uns_a / uns_b; $display("%1d",uns_r);
      $finish();
   end

endmodule
